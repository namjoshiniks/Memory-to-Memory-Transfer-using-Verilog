module Comparator_tb();

wire Sign;
reg [7:0] DOut1,DOut2;
reg clk;
 
always
#5 clk = ~clk;

Comparator MUT(DOut2,DOut1,Sign);

initial begin
clk = 1'b0;
DOut2 = 8'b00000000;
DOut1 = 8'b00000000;

@(posedge clk)
begin
 DOut2 = 8'b00000011;
 DOut1 = 8'b00000001;
end

@(posedge clk)
begin
 DOut2 = 8'b10000000;
 DOut1 = 8'b10000011;
end

@(posedge clk)
begin
 DOut2 = 8'b00000111;
 DOut1 = 8'b00010000;
end

@(posedge clk)
begin
 DOut2 = 8'b10011111;
 DOut1 = 8'b10001111;
end

@(posedge clk)
begin
 DOut2 = 8'b10000001;
 DOut1 = 8'b10000010;
end

end

endmodule